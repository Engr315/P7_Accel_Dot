`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
// Created for Indiana University's E315 Class
//
// 
// Andrew Lukefahr
// lukefahr@iu.edu
//
// 2021-03-24
//
//////////////////////////////////////////////////////////////////////////////////


module accel_dot_20_10_tb();

    integer                     i;
    
    // Clock signal
    bit                         clk;
    // Reset signal
    bit                         rst;

    // Incomming Matrix AXI4-Stream
    reg [31:0]                  INPUT_AXIS_TDATA;
    reg                         INPUT_AXIS_TLAST;
    reg                         INPUT_AXIS_TVALID;
    wire                        INPUT_AXIS_TREADY;
    
    // Outgoing Vector AXI4-Stream 		
    wire [31:0]                 OUTPUT_AXIS_TDATA;
    wire                        OUTPUT_AXIS_TLAST;
    wire                        OUTPUT_AXIS_TVALID;
    logic                       OUTPUT_AXIS_TREADY;

    // This is autogenerated. see python/dot_20_10.py for details. 
    localparam ROWS = 20;
    localparam COLS = 10;

    localparam logic [31:0] weights [0:ROWS-1] [0:COLS-1] = '{
      '{
        $shortrealtobits(0.025832674),$shortrealtobits(0.031067913),$shortrealtobits(0.074954145),$shortrealtobits(0.069431275),
        $shortrealtobits(0.027941115),$shortrealtobits(-0.38890076),$shortrealtobits(0.033413205),$shortrealtobits(0.023418507),
        $shortrealtobits(0.06414384),$shortrealtobits(0.03908126)
      },
      '{
        $shortrealtobits(0.47429913),$shortrealtobits(-0.030727461),$shortrealtobits(-0.07559153),$shortrealtobits(-0.06562075),
        $shortrealtobits(-0.027017677),$shortrealtobits(-0.1192499),$shortrealtobits(-0.033655476),$shortrealtobits(-0.023151854),
        $shortrealtobits(-0.06256888),$shortrealtobits(-0.038519256)
      },
      '{
        $shortrealtobits(0.11026208),$shortrealtobits(-0.21939886),$shortrealtobits(0.13531552),$shortrealtobits(0.032739077),
        $shortrealtobits(-0.100836486),$shortrealtobits(0.0315356),$shortrealtobits(-0.070727594),$shortrealtobits(-0.060791247),
        $shortrealtobits(0.109173514),$shortrealtobits(-0.09761812)
      },
      '{
        $shortrealtobits(-0.09525199),$shortrealtobits(-0.015320993),$shortrealtobits(0.27705696),$shortrealtobits(0.29808667),
        $shortrealtobits(-0.0757019),$shortrealtobits(-0.35671774),$shortrealtobits(-0.36361465),$shortrealtobits(-0.19701016),
        $shortrealtobits(0.07038336),$shortrealtobits(-0.065721996)
      },
      '{
        $shortrealtobits(-0.0054014125),$shortrealtobits(-0.0017534702),$shortrealtobits(-0.02180146),$shortrealtobits(-0.043511778),
        $shortrealtobits(0.0126061505),$shortrealtobits(-0.06802737),$shortrealtobits(-0.022320164),$shortrealtobits(0.05773446),
        $shortrealtobits(0.0007781352),$shortrealtobits(0.093098156)
      },
      '{
        $shortrealtobits(0.15577213),$shortrealtobits(0.34477082),$shortrealtobits(0.090137675),$shortrealtobits(-0.31324303),
        $shortrealtobits(-0.3665532),$shortrealtobits(0.020112142),$shortrealtobits(-0.17536488),$shortrealtobits(0.30936924),
        $shortrealtobits(-0.33058545),$shortrealtobits(-0.14599612)
      },
      '{
        $shortrealtobits(0.0833357),$shortrealtobits(0.35463968),$shortrealtobits(0.034455944),$shortrealtobits(-0.17448412),
        $shortrealtobits(-0.14407434),$shortrealtobits(0.34011856),$shortrealtobits(-0.37385958),$shortrealtobits(0.21625571),
        $shortrealtobits(-0.31103995),$shortrealtobits(0.045323063)
      },
      '{
        $shortrealtobits(-0.02596514),$shortrealtobits(-0.034139764),$shortrealtobits(-0.074281424),$shortrealtobits(-0.06537479),
        $shortrealtobits(-0.027002666),$shortrealtobits(-0.12030753),$shortrealtobits(-0.032794163),$shortrealtobits(-0.022686793),
        $shortrealtobits(0.443038),$shortrealtobits(-0.04100036)
      },
      '{
        $shortrealtobits(-0.020247536),$shortrealtobits(-0.028367976),$shortrealtobits(-0.05547012),$shortrealtobits(-0.02299753),
        $shortrealtobits(0.4642982),$shortrealtobits(-0.049594223),$shortrealtobits(-0.012405541),$shortrealtobits(-0.08192114),
        $shortrealtobits(-0.063603744),$shortrealtobits(-0.13136235)
      },
      '{
        $shortrealtobits(-0.08965313),$shortrealtobits(-0.015638348),$shortrealtobits(0.31165576),$shortrealtobits(-0.0017556128),
        $shortrealtobits(0.22123784),$shortrealtobits(-0.29498687),$shortrealtobits(0.12892826),$shortrealtobits(-0.059905306),
        $shortrealtobits(-0.26068124),$shortrealtobits(-0.14420311)
      },
      '{
        $shortrealtobits(-0.021710042),$shortrealtobits(-0.029718418),$shortrealtobits(-0.05677786),$shortrealtobits(-0.024768198),
        $shortrealtobits(-0.037383515),$shortrealtobits(-0.052242942),$shortrealtobits(-0.0105619235),$shortrealtobits(0.42426327),
        $shortrealtobits(-0.062348627),$shortrealtobits(-0.12969314)
      },
      '{
        $shortrealtobits(-0.33830196),$shortrealtobits(-0.21303433),$shortrealtobits(-0.048951115),$shortrealtobits(0.25440967),
        $shortrealtobits(-0.22557631),$shortrealtobits(-0.09242142),$shortrealtobits(-0.055013154),$shortrealtobits(0.37846345),
        $shortrealtobits(0.2120045),$shortrealtobits(-0.2063289)
      },
      '{
        $shortrealtobits(-0.0014902132),$shortrealtobits(-0.5039727),$shortrealtobits(0.508414),$shortrealtobits(-0.001196809),
        $shortrealtobits(0.00043627736),$shortrealtobits(-0.0005926093),$shortrealtobits(-0.0012271563),$shortrealtobits(-0.00072608533),
        $shortrealtobits(-0.000416694),$shortrealtobits(2.0524347e-05)
      },
      '{
        $shortrealtobits(-0.026448617),$shortrealtobits(-0.031083299),$shortrealtobits(-0.07606366),$shortrealtobits(0.43673903),
        $shortrealtobits(-0.026514161),$shortrealtobits(-0.11752776),$shortrealtobits(-0.032170594),$shortrealtobits(-0.022210078),
        $shortrealtobits(-0.06506433),$shortrealtobits(-0.03911492)
      },
      '{
        $shortrealtobits(0.35377282),$shortrealtobits(-0.3778204),$shortrealtobits(0.29622322),$shortrealtobits(0.02397883),
        $shortrealtobits(-0.3820959),$shortrealtobits(-0.223997),$shortrealtobits(-0.16420537),$shortrealtobits(0.10098358),
        $shortrealtobits(-0.056816496),$shortrealtobits(-0.11162076)
      },
      '{
        $shortrealtobits(0.020578936),$shortrealtobits(0.028920183),$shortrealtobits(0.05403632),$shortrealtobits(0.023214692),
        $shortrealtobits(0.041436687),$shortrealtobits(0.049547866),$shortrealtobits(0.01047655),$shortrealtobits(0.0813296),
        $shortrealtobits(0.0643888),$shortrealtobits(-0.3736555)
      },
      '{
        $shortrealtobits(-0.02662784),$shortrealtobits(-0.03034657),$shortrealtobits(-0.0781744),$shortrealtobits(-0.06629315),
        $shortrealtobits(-0.027823025),$shortrealtobits(-0.11695455),$shortrealtobits(0.46898773),$shortrealtobits(-0.021602403),
        $shortrealtobits(-0.06392121),$shortrealtobits(-0.038148273)
      },
      '{
        $shortrealtobits(-0.21310297),$shortrealtobits(0.200328),$shortrealtobits(-0.2060856),$shortrealtobits(-0.25261205),
        $shortrealtobits(-0.13819245),$shortrealtobits(0.01940004),$shortrealtobits(0.019376138),$shortrealtobits(0.2770613),
        $shortrealtobits(-0.33503842),$shortrealtobits(-0.13916487)
      },
      '{
        $shortrealtobits(0.38198224),$shortrealtobits(-0.24366285),$shortrealtobits(0.120944664),$shortrealtobits(0.01898678),
        $shortrealtobits(0.20554696),$shortrealtobits(0.040481124),$shortrealtobits(0.23627168),$shortrealtobits(-0.28644764),
        $shortrealtobits(0.22857712),$shortrealtobits(0.4494442)
      },
      '{
        $shortrealtobits(-0.028221987),$shortrealtobits(-0.033350915),$shortrealtobits(0.43056083),$shortrealtobits(-0.06829891),
        $shortrealtobits(-0.02646765),$shortrealtobits(-0.117585674),$shortrealtobits(-0.03333983),$shortrealtobits(-0.022141851),
        $shortrealtobits(-0.06445468),$shortrealtobits(-0.037462544)
        }
    };

    //used to access the FP tests table    
    bit [31:0] fp_hex;
    //used to access the FP Solutions table
    bit [31:0] sol_hex;
 
    reg COMPUTE_FIN;

    accel_dot #(
        .ROWS(ROWS),
        .COLS(COLS)
    ) DUT ( 
        .clk, 
        .rst, 

        .weights(weights),

        .INPUT_AXIS_TDATA,
        .INPUT_AXIS_TLAST,
        .INPUT_AXIS_TVALID,
        .INPUT_AXIS_TREADY,
        
        .OUTPUT_AXIS_TDATA,
        .OUTPUT_AXIS_TLAST,
        .OUTPUT_AXIS_TVALID,
        .OUTPUT_AXIS_TREADY

    );  


    always #10 clk <= ~clk;
    
    // see python/dot_20_10.py for values
    task inputs_table_lookup(
        input integer id,
        output bit [31:0] hex
        );

        static bit [31:0] fpHex [0:19] = {
         $shortrealtobits(0.9992157677176247), $shortrealtobits(-0.9992391649984632), $shortrealtobits(-0.996713106729648),
         $shortrealtobits(-0.9989178474188565), $shortrealtobits(-0.9991897304310112), $shortrealtobits(-0.9992238976312111),
         $shortrealtobits(-0.999874794745124), $shortrealtobits(-0.9999983469326711), $shortrealtobits(-0.9999823366958234),
         $shortrealtobits(-0.9993464993540697), $shortrealtobits(-0.99999895931321), $shortrealtobits(-0.9994030383922219),
         $shortrealtobits(0.999932362106602), $shortrealtobits(-0.9999615682027578), $shortrealtobits(0.9981479711735248),
         $shortrealtobits(0.9997359101642), $shortrealtobits(0.9966997506542944), $shortrealtobits(0.9973577360650924),
         $shortrealtobits(-0.9991081374552344), $shortrealtobits(-0.9924563156913059)
        };
        static int MAX_SIZE = 20;

        assert(id < MAX_SIZE) else $fatal(1, "Bad id");
        hex = fpHex[id];
    endtask : inputs_table_lookup  
    
    // see python/dot_20_10.py for values
    task outputs_table_lookup(
        input integer id,
        output bit [31:0] hex
        );

        static bit [31:0] fpHex [0:9] = {
         $shortrealtobits(-0.39490294817324495), $shortrealtobits(-0.4558233633141949), $shortrealtobits(-0.3374061380803292),
         $shortrealtobits(-0.463853652749869), $shortrealtobits(-0.3244523604970557), $shortrealtobits(0.29448396778040775),
         $shortrealtobits(1.215281511185426), $shortrealtobits(-0.1505974181548544), $shortrealtobits(-0.17037033565393786),
         $shortrealtobits(-0.1341205480148839)
        };
        static int MAX_SIZE = 10;

                
        assert(id <MAX_SIZE) else $fatal(1, "Bad id");
        hex = fpHex[id];
    endtask: outputs_table_lookup
    
    
    task send_word_axi4stream(
        input logic [31:0] data,
        input logic last
    );
    
        INPUT_AXIS_TDATA = data;
        INPUT_AXIS_TVALID='h1;
        INPUT_AXIS_TLAST = last;
        #1;
        while( INPUT_AXIS_TREADY == 'h0)  begin
            @(negedge clk);
            #1;
        end
        
        @(negedge clk);
        INPUT_AXIS_TVALID='h0;
        INPUT_AXIS_TLAST='h0;

    endtask

    task recv_word_axi4stream(
        output logic [31:0] data
    );
    
        OUTPUT_AXIS_TREADY = 'h1;
        #1;
        while (OUTPUT_AXIS_TVALID == 'h0) begin
            @(negedge clk);
            #1;
        end
        
        data = OUTPUT_AXIS_TDATA;
        @(negedge clk);
        OUTPUT_AXIS_TREADY = 'h0;
    
    endtask    

    task init();

        clk = 'h0;
        rst = 'h1;

        INPUT_AXIS_TDATA = 'h0;
        INPUT_AXIS_TLAST = 'h0;
        INPUT_AXIS_TVALID = 'h0;
        
        OUTPUT_AXIS_TREADY = 'h0;
      
       i = 0;
    endtask

    task compute();
         
        COMPUTE_FIN = 'h0;

        $display("Sending Input Vector");                
        for (i = 0; i < ROWS; ++i) begin
            inputs_table_lookup(i, fp_hex);
            $display( "Sending %h (%f)", fp_hex, $bitstoshortreal(fp_hex) ); 
            send_word_axi4stream(fp_hex, i == 19);
        end                
              
        $display("Receiving Output Vector");
        for (i = 0; i < COLS; ++i) begin
            real mismatch; 
            
            outputs_table_lookup(i, sol_hex);
            
            recv_word_axi4stream(fp_hex);
            
            $display( "Received %h (%f)",
                fp_hex, $bitstoshortreal(fp_hex));
             //compute the difference between what was observed and what was
            // expected with Python
            mismatch = $bitstoshortreal(fp_hex) - $bitstoshortreal(sol_hex);
            $display("mismatch: %f", mismatch);
            
            assert( (mismatch > -0.000001) && (mismatch < +0.000001) ) else
                $fatal(1, "Bad Test Response %h (%f), Expected %h (%f) mismatch:%f", 
                    fp_hex, $bitstoshortreal(fp_hex), sol_hex, $bitstoshortreal(sol_hex), mismatch); 
    
            //pause the output stream after each value            
            OUTPUT_AXIS_TREADY='h0;
            repeat(2) @(negedge clk);

        end
        $display( "Compute done, finish timing" );
        COMPUTE_FIN = 'h1;
    endtask

    task timeit (
        output int cycles
        );
        
        cycles = 0;
        while ( ! (
            (OUTPUT_AXIS_TREADY === 'h1) && 
            (OUTPUT_AXIS_TVALID === 'h1) && 
            (OUTPUT_AXIS_TLAST === 'h1) ) ) begin
            cycles += 1;
            
            @(posedge clk);
            
            assert (cycles < 44100) else 
                $fatal(1, "Running too long, check OUTPUT_AXIS?");
        end
                        
        @(posedge clk);
        assert(COMPUTE_FIN == 'h1) else
            $fatal(1, "Timing done before correctness check");

    endtask
    

    //Main process
    initial begin
 
        int cycles;
        
        $timeformat (-12, 1, " ps", 1);      

        $display("Simulation Setup");
        init();
        
        $display("Holding Reset");
        for (i = 0; i < 20; i++) 
        @(negedge clk);

        rst = 0;        

        repeat(2) @(negedge clk);
        
        $display("Starting Simulation");
        $display("NOTE:  this one has extra delays"); 
        
        fork
            compute();
            timeit(cycles);
        join                                                  
        
        $display("@@@Passed in %d Cycles (was 2210)", cycles);
        
        $finish;

    end

endmodule
